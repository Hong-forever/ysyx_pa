module scpu
(

);


endmodule
