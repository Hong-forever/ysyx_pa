module top
#(
    parameter DATA_WIDTH = 8
)(
    input   wire                  clk,
    input   wire                  rstn,
    
    input   wire                  ps2_clk,
    input   wire                  ps2_data,
    
    output  wire                  ready,
    output  wire                  overflow,
    
    output  wire [7:0]            seg0,
    output  wire [7:0]            seg1,
    output  wire [7:0]            seg2,
    output  wire [7:0]            seg3,
    output  wire [7:0]            seg4,
    output  wire [7:0]            seg5,
    output  wire [7:0]            seg6,
    output  wire [7:0]            seg7
);

    wire [7:0] key_code;
    reg [7:0] ascii;
    reg next_data;
    
    always @(posedge clk) begin
        if(rstn) next_data <= 1'b1;
        else if(ready) next_data <= 1'b0;
        else next_data <= 1'b1;
    end

    ps2_key ps2_key_inst
    (
        .clk                (clk        ),
        .clrn               (rstn       ),
        .ps2_clk            (ps2_clk    ),
        .ps2_data           (ps2_data   ),
        .data               (key_code   ),
        .ready              (ready      ),
        .nextdata_n         (next_data  ),
        .overflow           (overflow   )
    );
    
    always @(*) begin
        case(key_code)
            8'h45: ascii = 8'h30; // 0
            8'h16: ascii = 8'h31; // 1
            8'h1E: ascii = 8'h32; // 2
            8'h26: ascii = 8'h33; // 3
            8'h25: ascii = 8'h34; // 4
            8'h2E: ascii = 8'h35; // 5
            8'h36: ascii = 8'h36; // 6
            8'h3D: ascii = 8'h37; // 7
            8'h3E: ascii = 8'h38; // 8
            8'h46: ascii = 8'h39; // 9
        
            // 小写字母 a-z
            8'h1C: ascii = 8'h61; // a
            8'h32: ascii = 8'h62; // b
            8'h21: ascii = 8'h63; // c
            8'h23: ascii = 8'h64; // d
            8'h24: ascii = 8'h65; // e
            8'h2B: ascii = 8'h66; // f
            8'h34: ascii = 8'h67; // g
            8'h33: ascii = 8'h68; // h
            8'h43: ascii = 8'h69; // i
            8'h3B: ascii = 8'h6A; // j
            8'h42: ascii = 8'h6B; // k
            8'h4B: ascii = 8'h6C; // l
            8'h3A: ascii = 8'h6D; // m
            8'h31: ascii = 8'h6E; // n
            8'h44: ascii = 8'h6F; // o
            8'h4D: ascii = 8'h70; // p
            8'h15: ascii = 8'h71; // q
            8'h2D: ascii = 8'h72; // r
            8'h1B: ascii = 8'h73; // s
            8'h2C: ascii = 8'h74; // t
            8'h3C: ascii = 8'h75; // u
            8'h2A: ascii = 8'h76; // v
            8'h1D: ascii = 8'h77; // w
            8'h22: ascii = 8'h78; // x
            8'h35: ascii = 8'h79; // y
            8'h1A: ascii = 8'h7A; // z
            default: ascii = 8'hff;
        endcase
    end
    
    

    segs segs_inst0
    (
        .din                (key_code   ),

        .seg0               (seg0       ),
        .seg1               (seg1       )
    );
    
    segs segs_inst1
    (
        .din                (ascii      ),

        .seg0               (seg2       ),
        .seg1               (seg3       )
    );
    
    segs segs_inst2
    (
        .din                (0   ),

        .seg0               (seg4       ),
        .seg1               (seg5       )
    );
    
    segs segs_inst3
    (
        .din                (0   ),

        .seg0               (seg6       ),
        .seg1               (seg7       )
    );
    
endmodule
